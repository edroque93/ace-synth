module mem_stage (
);
endmodule
