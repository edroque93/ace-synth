module id_stage (
);
endmodule
