module ex_stage (
);
endmodule
